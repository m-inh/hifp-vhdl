library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.dwt_pkg.all;

entity hifp_tb is
    generic (num_of_fpid_frames : positive := 2);
end entity;

architecture rtl of hifp_tb is

    signal tb_wave_all: natural_array(0 to num_of_fpid_frames*32-1);
    signal tb_fpid_all: std_logic_vector(0 to num_of_fpid_frames-1);

    component hifp is
        generic (num_of_fpid_frames: positive);
    
        port (
            wave_all: in natural_array(0 to num_of_fpid_frames*32-1);
            fpid_all: out std_logic_vector(0 to num_of_fpid_frames-1)
        );
    end component;

begin

    en_hifp: hifp
    generic map (num_of_fpid_frames => num_of_fpid_frames)
    port map (
        tb_wave_all,
        tb_fpid_all
    );

    process is
    begin
        -- tb_wave_all <= (1, 1, 1, 1, 1, 1, 1, 1, others => 0);
        -- wait for 100 ns;

        -- tb_wave_all(0) <= 3;
        -- tb_wave_all(1) <= 3;
        -- tb_wave_all(2) <= 3;
        -- tb_wave_all(3) <= 3;
        -- tb_wave_all(4) <= 3;
        -- tb_wave_all(5) <= 3;
        -- tb_wave_all(6) <= 3;
        -- tb_wave_all(7) <= 3;
        -- tb_wave_all(8) <= 2;
        -- tb_wave_all(9) <= 2;
        -- tb_wave_all(10) <= 2;
        -- tb_wave_all(11) <= 2;
        -- tb_wave_all(12) <= 2;
        -- tb_wave_all(13) <= 2;
        -- tb_wave_all(14) <= 2;
        -- tb_wave_all(15) <= 2;
        -- tb_wave_all(16) <= 2;
        -- tb_wave_all(17) <= 2;
        -- tb_wave_all(18) <= 2;
        -- tb_wave_all(19) <= 2;
        -- tb_wave_all(20) <= 2;
        -- tb_wave_all(21) <= 2;
        -- tb_wave_all(22) <= 2;
        -- tb_wave_all(23) <= 2;
        -- tb_wave_all(24) <= 2;
        -- tb_wave_all(25) <= 2;
        -- tb_wave_all(26) <= 2;
        -- tb_wave_all(27) <= 2;
        -- tb_wave_all(28) <= 2;
        -- tb_wave_all(29) <= 2;
        -- tb_wave_all(30) <= 2;
        -- tb_wave_all(31) <= 2;

        -- tb_wave_all(32) <= 4;
        -- tb_wave_all(33) <= 4;
        -- tb_wave_all(34) <= 4;
        -- tb_wave_all(35) <= 4;
        -- tb_wave_all(36) <= 4;
        -- tb_wave_all(37) <= 4;
        -- tb_wave_all(38) <= 4;
        -- tb_wave_all(39) <= 4;
        -- tb_wave_all(40) <= 2;
        -- tb_wave_all(41) <= 2;
        -- tb_wave_all(42) <= 2;
        -- tb_wave_all(43) <= 2;
        -- tb_wave_all(44) <= 2;
        -- tb_wave_all(45) <= 2;
        -- tb_wave_all(46) <= 2;
        -- tb_wave_all(47) <= 2;
        -- tb_wave_all(48) <= 2;
        -- tb_wave_all(49) <= 2;
        -- tb_wave_all(50) <= 2;
        -- tb_wave_all(51) <= 2;
        -- tb_wave_all(52) <= 2;
        -- tb_wave_all(53) <= 2;
        -- tb_wave_all(54) <= 2;
        -- tb_wave_all(55) <= 2;
        -- tb_wave_all(56) <= 2;
        -- tb_wave_all(57) <= 2;
        -- tb_wave_all(58) <= 2;
        -- tb_wave_all(59) <= 2;
        -- tb_wave_all(60) <= 2;
        -- tb_wave_all(61) <= 2;
        -- tb_wave_all(62) <= 2;
        -- tb_wave_all(63) <= 2;
        
        -- wait for 100 ns;
        

        -- tb_wave_all <= (1, 2, 3, 4, 5, 6, 7, 8, others => 7);
        -- wait for 100 ns;



        tb_wave_all(0) <= 0; 
        tb_wave_all(1) <= 0; 
        tb_wave_all(2) <= 0; 
        tb_wave_all(3) <= 0; 
        tb_wave_all(4) <= 0; 
        tb_wave_all(5) <= 0; 
        tb_wave_all(6) <= 0; 
        tb_wave_all(7) <= 0; 
        tb_wave_all(8) <= 0; 
        tb_wave_all(9) <= 0; 
        tb_wave_all(10) <= 0; 
        tb_wave_all(11) <= 0; 
        tb_wave_all(12) <= 0; 
        tb_wave_all(13) <= 0; 
        tb_wave_all(14) <= 0; 
        tb_wave_all(15) <= 0; 
        tb_wave_all(16) <= 0; 
        tb_wave_all(17) <= 0; 
        tb_wave_all(18) <= 0; 
        tb_wave_all(19) <= 0; 
        tb_wave_all(20) <= 0; 
        tb_wave_all(21) <= 0; 
        tb_wave_all(22) <= 0; 
        tb_wave_all(23) <= 0; 
        tb_wave_all(24) <= 0; 
        tb_wave_all(25) <= 0; 
        tb_wave_all(26) <= 0; 
        tb_wave_all(27) <= 0; 
        tb_wave_all(28) <= 0; 
        tb_wave_all(29) <= 0; 
        tb_wave_all(30) <= 0; 
        tb_wave_all(31) <= 0; 
        tb_wave_all(32) <= 0; 
        tb_wave_all(33) <= 0; 
        tb_wave_all(34) <= 0; 
        tb_wave_all(35) <= 0; 
        tb_wave_all(36) <= 0; 
        tb_wave_all(37) <= 0; 
        tb_wave_all(38) <= 0; 
        tb_wave_all(39) <= 0; 
        tb_wave_all(40) <= 0; 
        tb_wave_all(41) <= 0; 
        tb_wave_all(42) <= 0; 
        tb_wave_all(43) <= 0; 
        tb_wave_all(44) <= 0; 
        tb_wave_all(45) <= 0; 
        tb_wave_all(46) <= 0; 
        tb_wave_all(47) <= 0; 
        tb_wave_all(48) <= 0; 
        tb_wave_all(49) <= 0; 
        tb_wave_all(50) <= 0; 
        tb_wave_all(51) <= 0; 
        tb_wave_all(52) <= 0; 
        tb_wave_all(53) <= 0; 
        tb_wave_all(54) <= 0; 
        tb_wave_all(55) <= 0; 
        tb_wave_all(56) <= 0; 
        tb_wave_all(57) <= 0; 
        tb_wave_all(58) <= 0; 
        tb_wave_all(59) <= 0; 
        tb_wave_all(60) <= 0; 
        tb_wave_all(61) <= 0; 
        tb_wave_all(62) <= 0; 
        tb_wave_all(63) <= 0; 
        tb_wave_all(64) <= 0; 
        tb_wave_all(65) <= 65533; 
        tb_wave_all(66) <= 7; 
        tb_wave_all(67) <= 3; 
        tb_wave_all(68) <= 65518; 
        tb_wave_all(69) <= 9; 
        tb_wave_all(70) <= 65532; 
        tb_wave_all(71) <= 65497; 
        tb_wave_all(72) <= 0; 
        tb_wave_all(73) <= 0; 
        tb_wave_all(74) <= 0; 
        tb_wave_all(75) <= 0; 
        tb_wave_all(76) <= 0; 
        tb_wave_all(77) <= 0; 
        tb_wave_all(78) <= 0; 
        tb_wave_all(79) <= 0; 
        tb_wave_all(80) <= 0; 
        tb_wave_all(81) <= 0; 
        tb_wave_all(82) <= 0; 
        tb_wave_all(83) <= 0; 
        tb_wave_all(84) <= 0; 
        tb_wave_all(85) <= 0; 
        tb_wave_all(86) <= 0; 
        tb_wave_all(87) <= 0; 
        tb_wave_all(88) <= 0; 
        tb_wave_all(89) <= 0; 
        tb_wave_all(90) <= 0; 
        tb_wave_all(91) <= 0; 
        tb_wave_all(92) <= 0; 
        tb_wave_all(93) <= 0; 
        tb_wave_all(94) <= 0; 
        tb_wave_all(95) <= 0; 
        tb_wave_all(96) <= 1591; 
        tb_wave_all(97) <= 1586; 
        tb_wave_all(98) <= 1999; 
        tb_wave_all(99) <= 1963; 
        tb_wave_all(100) <= 1521; 
        tb_wave_all(101) <= 1130; 
        tb_wave_all(102) <= 1204; 
        tb_wave_all(103) <= 718; 
        tb_wave_all(104) <= 0; 
        tb_wave_all(105) <= 0; 
        tb_wave_all(106) <= 0; 
        tb_wave_all(107) <= 0; 
        tb_wave_all(108) <= 0; 
        tb_wave_all(109) <= 0; 
        tb_wave_all(110) <= 0; 
        tb_wave_all(111) <= 0; 
        tb_wave_all(112) <= 0; 
        tb_wave_all(113) <= 0; 
        tb_wave_all(114) <= 0; 
        tb_wave_all(115) <= 0; 
        tb_wave_all(116) <= 0; 
        tb_wave_all(117) <= 0; 
        tb_wave_all(118) <= 0; 
        tb_wave_all(119) <= 0; 
        tb_wave_all(120) <= 0; 
        tb_wave_all(121) <= 0; 
        tb_wave_all(122) <= 0; 
        tb_wave_all(123) <= 0; 
        tb_wave_all(124) <= 0; 
        tb_wave_all(125) <= 0; 
        tb_wave_all(126) <= 0; 
        tb_wave_all(127) <= 0; 
        tb_wave_all(128) <= 63660; 
        tb_wave_all(129) <= 63902; 
        tb_wave_all(130) <= 64374; 
        tb_wave_all(131) <= 64602; 
        tb_wave_all(132) <= 65070; 
        tb_wave_all(133) <= 65264; 
        tb_wave_all(134) <= 65145; 
        tb_wave_all(135) <= 65496; 
        tb_wave_all(136) <= 0; 
        tb_wave_all(137) <= 0; 
        tb_wave_all(138) <= 0; 
        tb_wave_all(139) <= 0; 
        tb_wave_all(140) <= 0; 
        tb_wave_all(141) <= 0; 
        tb_wave_all(142) <= 0; 
        tb_wave_all(143) <= 0; 
        tb_wave_all(144) <= 0; 
        tb_wave_all(145) <= 0; 
        tb_wave_all(146) <= 0; 
        tb_wave_all(147) <= 0; 
        tb_wave_all(148) <= 0; 
        tb_wave_all(149) <= 0; 
        tb_wave_all(150) <= 0; 
        tb_wave_all(151) <= 0; 
        tb_wave_all(152) <= 0; 
        tb_wave_all(153) <= 0; 
        tb_wave_all(154) <= 0; 
        tb_wave_all(155) <= 0; 
        tb_wave_all(156) <= 0; 
        tb_wave_all(157) <= 0; 
        tb_wave_all(158) <= 0; 
        tb_wave_all(159) <= 0; 
        tb_wave_all(160) <= 1079; 
        tb_wave_all(161) <= 1815; 
        tb_wave_all(162) <= 1818; 
        tb_wave_all(163) <= 985; 
        tb_wave_all(164) <= 999; 
        tb_wave_all(165) <= 1284; 
        tb_wave_all(166) <= 1634; 
        tb_wave_all(167) <= 1419; 
        tb_wave_all(168) <= 0; 
        tb_wave_all(169) <= 0; 
        tb_wave_all(170) <= 0; 
        tb_wave_all(171) <= 0; 
        tb_wave_all(172) <= 0; 
        tb_wave_all(173) <= 0; 
        tb_wave_all(174) <= 0; 
        tb_wave_all(175) <= 0; 
        tb_wave_all(176) <= 0; 
        tb_wave_all(177) <= 0; 
        tb_wave_all(178) <= 0; 
        tb_wave_all(179) <= 0; 
        tb_wave_all(180) <= 0; 
        tb_wave_all(181) <= 0; 
        tb_wave_all(182) <= 0; 
        tb_wave_all(183) <= 0; 
        tb_wave_all(184) <= 0; 
        tb_wave_all(185) <= 0; 
        tb_wave_all(186) <= 0; 
        tb_wave_all(187) <= 0; 
        tb_wave_all(188) <= 0; 
        tb_wave_all(189) <= 0; 
        tb_wave_all(190) <= 0; 
        tb_wave_all(191) <= 0; 
        tb_wave_all(192) <= 2981; 
        tb_wave_all(193) <= 2882; 
        tb_wave_all(194) <= 1504; 
        tb_wave_all(195) <= 1095; 
        tb_wave_all(196) <= 1452; 
        tb_wave_all(197) <= 1579; 
        tb_wave_all(198) <= 1452; 
        tb_wave_all(199) <= 544; 
        tb_wave_all(200) <= 0; 
        tb_wave_all(201) <= 0; 
        tb_wave_all(202) <= 0; 
        tb_wave_all(203) <= 0; 
        tb_wave_all(204) <= 0; 
        tb_wave_all(205) <= 0; 
        tb_wave_all(206) <= 0; 
        tb_wave_all(207) <= 0; 
        tb_wave_all(208) <= 0; 
        tb_wave_all(209) <= 0; 
        tb_wave_all(210) <= 0; 
        tb_wave_all(211) <= 0; 
        tb_wave_all(212) <= 0; 
        tb_wave_all(213) <= 0; 
        tb_wave_all(214) <= 0; 
        tb_wave_all(215) <= 0; 
        tb_wave_all(216) <= 0; 
        tb_wave_all(217) <= 0; 
        tb_wave_all(218) <= 0; 
        tb_wave_all(219) <= 0; 
        tb_wave_all(220) <= 0; 
        tb_wave_all(221) <= 0; 
        tb_wave_all(222) <= 0; 
        tb_wave_all(223) <= 0; 
        tb_wave_all(224) <= 63764; 
        tb_wave_all(225) <= 63942; 
        tb_wave_all(226) <= 62380; 
        tb_wave_all(227) <= 63195; 
        tb_wave_all(228) <= 63409; 
        tb_wave_all(229) <= 62323; 
        tb_wave_all(230) <= 62649; 
        tb_wave_all(231) <= 63559; 
        tb_wave_all(232) <= 0; 
        tb_wave_all(233) <= 0; 
        tb_wave_all(234) <= 0; 
        tb_wave_all(235) <= 0; 
        tb_wave_all(236) <= 0; 
        tb_wave_all(237) <= 0; 
        tb_wave_all(238) <= 0; 
        tb_wave_all(239) <= 0; 
        tb_wave_all(240) <= 0; 
        tb_wave_all(241) <= 0; 
        tb_wave_all(242) <= 0; 
        tb_wave_all(243) <= 0; 
        tb_wave_all(244) <= 0; 
        tb_wave_all(245) <= 0; 
        tb_wave_all(246) <= 0; 
        tb_wave_all(247) <= 0; 
        tb_wave_all(248) <= 0; 
        tb_wave_all(249) <= 0; 
        tb_wave_all(250) <= 0; 
        tb_wave_all(251) <= 0; 
        tb_wave_all(252) <= 0; 
        tb_wave_all(253) <= 0; 
        tb_wave_all(254) <= 0; 
        tb_wave_all(255) <= 0; 
        tb_wave_all(256) <= 36; 
        tb_wave_all(257) <= 773; 
        tb_wave_all(258) <= 1131; 
        tb_wave_all(259) <= 758; 
        tb_wave_all(260) <= 737; 
        tb_wave_all(261) <= 1465; 
        tb_wave_all(262) <= 1486; 
        tb_wave_all(263) <= 762; 
        tb_wave_all(264) <= 0; 
        tb_wave_all(265) <= 0; 
        tb_wave_all(266) <= 0; 
        tb_wave_all(267) <= 0; 
        tb_wave_all(268) <= 0; 
        tb_wave_all(269) <= 0; 
        tb_wave_all(270) <= 0; 
        tb_wave_all(271) <= 0; 
        tb_wave_all(272) <= 0; 
        tb_wave_all(273) <= 0; 
        tb_wave_all(274) <= 0; 
        tb_wave_all(275) <= 0; 
        tb_wave_all(276) <= 0; 
        tb_wave_all(277) <= 0; 
        tb_wave_all(278) <= 0; 
        tb_wave_all(279) <= 0; 
        tb_wave_all(280) <= 0; 
        tb_wave_all(281) <= 0; 
        tb_wave_all(282) <= 0; 
        tb_wave_all(283) <= 0; 
        tb_wave_all(284) <= 0; 
        tb_wave_all(285) <= 0; 
        tb_wave_all(286) <= 0; 
        tb_wave_all(287) <= 0; 
        tb_wave_all(288) <= 302; 
        tb_wave_all(289) <= 228; 
        tb_wave_all(290) <= 2128; 
        tb_wave_all(291) <= 1855; 
        tb_wave_all(292) <= 2351; 
        tb_wave_all(293) <= 3377; 
        tb_wave_all(294) <= 2656; 
        tb_wave_all(295) <= 2260; 
        tb_wave_all(296) <= 0; 
        tb_wave_all(297) <= 0; 
        tb_wave_all(298) <= 0; 
        tb_wave_all(299) <= 0; 
        tb_wave_all(300) <= 0; 
        tb_wave_all(301) <= 0; 
        tb_wave_all(302) <= 0; 
        tb_wave_all(303) <= 0; 
        tb_wave_all(304) <= 0; 
        tb_wave_all(305) <= 0; 
        tb_wave_all(306) <= 0; 
        tb_wave_all(307) <= 0; 
        tb_wave_all(308) <= 0; 
        tb_wave_all(309) <= 0; 
        tb_wave_all(310) <= 0; 
        tb_wave_all(311) <= 0; 
        tb_wave_all(312) <= 0; 
        tb_wave_all(313) <= 0; 
        tb_wave_all(314) <= 0; 
        tb_wave_all(315) <= 0; 
        tb_wave_all(316) <= 0; 
        tb_wave_all(317) <= 0; 
        tb_wave_all(318) <= 0; 
        tb_wave_all(319) <= 0; 
        tb_wave_all(320) <= 65534; 
        tb_wave_all(321) <= 853; 
        tb_wave_all(322) <= 209; 
        tb_wave_all(323) <= 497; 
        tb_wave_all(324) <= 1738; 
        tb_wave_all(325) <= 725; 
        tb_wave_all(326) <= 65077; 
        tb_wave_all(327) <= 230; 
        tb_wave_all(328) <= 0; 
        tb_wave_all(329) <= 0; 
        tb_wave_all(330) <= 0; 
        tb_wave_all(331) <= 0; 
        tb_wave_all(332) <= 0; 
        tb_wave_all(333) <= 0; 
        tb_wave_all(334) <= 0; 
        tb_wave_all(335) <= 0; 
        tb_wave_all(336) <= 0; 
        tb_wave_all(337) <= 0; 
        tb_wave_all(338) <= 0; 
        tb_wave_all(339) <= 0; 
        tb_wave_all(340) <= 0; 
        tb_wave_all(341) <= 0; 
        tb_wave_all(342) <= 0; 
        tb_wave_all(343) <= 0; 
        tb_wave_all(344) <= 0; 
        tb_wave_all(345) <= 0; 
        tb_wave_all(346) <= 0; 
        tb_wave_all(347) <= 0; 
        tb_wave_all(348) <= 0; 
        tb_wave_all(349) <= 0; 
        tb_wave_all(350) <= 0; 
        tb_wave_all(351) <= 0; 
        tb_wave_all(352) <= 64067; 
        tb_wave_all(353) <= 63980; 
        tb_wave_all(354) <= 63076; 
        tb_wave_all(355) <= 65177; 
        tb_wave_all(356) <= 239; 
        tb_wave_all(357) <= 64424; 
        tb_wave_all(358) <= 64713; 
        tb_wave_all(359) <= 64635; 
        tb_wave_all(360) <= 0; 
        tb_wave_all(361) <= 0; 
        tb_wave_all(362) <= 0; 
        tb_wave_all(363) <= 0; 
        tb_wave_all(364) <= 0; 
        tb_wave_all(365) <= 0; 
        tb_wave_all(366) <= 0; 
        tb_wave_all(367) <= 0; 
        tb_wave_all(368) <= 0; 
        tb_wave_all(369) <= 0; 
        tb_wave_all(370) <= 0; 
        tb_wave_all(371) <= 0; 
        tb_wave_all(372) <= 0; 
        tb_wave_all(373) <= 0; 
        tb_wave_all(374) <= 0; 
        tb_wave_all(375) <= 0; 
        tb_wave_all(376) <= 0; 
        tb_wave_all(377) <= 0; 
        tb_wave_all(378) <= 0; 
        tb_wave_all(379) <= 0; 
        tb_wave_all(380) <= 0; 
        tb_wave_all(381) <= 0; 
        tb_wave_all(382) <= 0; 
        tb_wave_all(383) <= 0; 
        tb_wave_all(384) <= 1189; 
        tb_wave_all(385) <= 1168; 
        tb_wave_all(386) <= 430; 
        tb_wave_all(387) <= 688; 
        tb_wave_all(388) <= 1380; 
        tb_wave_all(389) <= 1023; 
        tb_wave_all(390) <= 1589; 
        tb_wave_all(391) <= 3386; 
        tb_wave_all(392) <= 0; 
        tb_wave_all(393) <= 0; 
        tb_wave_all(394) <= 0; 
        tb_wave_all(395) <= 0; 
        tb_wave_all(396) <= 0; 
        tb_wave_all(397) <= 0; 
        tb_wave_all(398) <= 0; 
        tb_wave_all(399) <= 0; 
        tb_wave_all(400) <= 0; 
        tb_wave_all(401) <= 0; 
        tb_wave_all(402) <= 0; 
        tb_wave_all(403) <= 0; 
        tb_wave_all(404) <= 0; 
        tb_wave_all(405) <= 0; 
        tb_wave_all(406) <= 0; 
        tb_wave_all(407) <= 0; 
        tb_wave_all(408) <= 0; 
        tb_wave_all(409) <= 0; 
        tb_wave_all(410) <= 0; 
        tb_wave_all(411) <= 0; 
        tb_wave_all(412) <= 0; 
        tb_wave_all(413) <= 0; 
        tb_wave_all(414) <= 0; 
        tb_wave_all(415) <= 0; 
        tb_wave_all(416) <= 63212; 
        tb_wave_all(417) <= 62089; 
        tb_wave_all(418) <= 62917; 
        tb_wave_all(419) <= 62813; 
        tb_wave_all(420) <= 62526; 
        tb_wave_all(421) <= 63789; 
        tb_wave_all(422) <= 63943; 
        tb_wave_all(423) <= 63757; 
        tb_wave_all(424) <= 0; 
        tb_wave_all(425) <= 0; 
        tb_wave_all(426) <= 0; 
        tb_wave_all(427) <= 0; 
        tb_wave_all(428) <= 0; 
        tb_wave_all(429) <= 0; 
        tb_wave_all(430) <= 0; 
        tb_wave_all(431) <= 0; 
        tb_wave_all(432) <= 0; 
        tb_wave_all(433) <= 0; 
        tb_wave_all(434) <= 0; 
        tb_wave_all(435) <= 0; 
        tb_wave_all(436) <= 0; 
        tb_wave_all(437) <= 0; 
        tb_wave_all(438) <= 0; 
        tb_wave_all(439) <= 0; 
        tb_wave_all(440) <= 0; 
        tb_wave_all(441) <= 0; 
        tb_wave_all(442) <= 0; 
        tb_wave_all(443) <= 0; 
        tb_wave_all(444) <= 0; 
        tb_wave_all(445) <= 0; 
        tb_wave_all(446) <= 0; 
        tb_wave_all(447) <= 0; 
        tb_wave_all(448) <= 171; 
        tb_wave_all(449) <= 65135; 
        tb_wave_all(450) <= 64304; 
        tb_wave_all(451) <= 64184; 
        tb_wave_all(452) <= 64859; 
        tb_wave_all(453) <= 64914; 
        tb_wave_all(454) <= 64599; 
        tb_wave_all(455) <= 63550; 
        tb_wave_all(456) <= 0; 
        tb_wave_all(457) <= 0; 
        tb_wave_all(458) <= 0; 
        tb_wave_all(459) <= 0; 
        tb_wave_all(460) <= 0; 
        tb_wave_all(461) <= 0; 
        tb_wave_all(462) <= 0; 
        tb_wave_all(463) <= 0; 
        tb_wave_all(464) <= 0; 
        tb_wave_all(465) <= 0; 
        tb_wave_all(466) <= 0; 
        tb_wave_all(467) <= 0; 
        tb_wave_all(468) <= 0; 
        tb_wave_all(469) <= 0; 
        tb_wave_all(470) <= 0; 
        tb_wave_all(471) <= 0; 
        tb_wave_all(472) <= 0; 
        tb_wave_all(473) <= 0; 
        tb_wave_all(474) <= 0; 
        tb_wave_all(475) <= 0; 
        tb_wave_all(476) <= 0; 
        tb_wave_all(477) <= 0; 
        tb_wave_all(478) <= 0; 
        tb_wave_all(479) <= 0; 
        tb_wave_all(480) <= 64352; 
        tb_wave_all(481) <= 356; 
        tb_wave_all(482) <= 838; 
        tb_wave_all(483) <= 65330; 
        tb_wave_all(484) <= 14; 
        tb_wave_all(485) <= 560; 
        tb_wave_all(486) <= 1147; 
        tb_wave_all(487) <= 942; 
        tb_wave_all(488) <= 0; 
        tb_wave_all(489) <= 0; 
        tb_wave_all(490) <= 0; 
        tb_wave_all(491) <= 0; 
        tb_wave_all(492) <= 0; 
        tb_wave_all(493) <= 0; 
        tb_wave_all(494) <= 0; 
        tb_wave_all(495) <= 0; 
        tb_wave_all(496) <= 0; 
        tb_wave_all(497) <= 0; 
        tb_wave_all(498) <= 0; 
        tb_wave_all(499) <= 0; 
        tb_wave_all(500) <= 0; 
        tb_wave_all(501) <= 0; 
        tb_wave_all(502) <= 0; 
        tb_wave_all(503) <= 0; 
        tb_wave_all(504) <= 0; 
        tb_wave_all(505) <= 0; 
        tb_wave_all(506) <= 0; 
        tb_wave_all(507) <= 0; 
        tb_wave_all(508) <= 0; 
        tb_wave_all(509) <= 0; 
        tb_wave_all(510) <= 0; 
        tb_wave_all(511) <= 0; 
        tb_wave_all(512) <= 63704; 
        tb_wave_all(513) <= 63661; 
        tb_wave_all(514) <= 63808; 
        tb_wave_all(515) <= 63573; 
        tb_wave_all(516) <= 63307; 
        tb_wave_all(517) <= 62858; 
        tb_wave_all(518) <= 62658; 
        tb_wave_all(519) <= 63579; 
        tb_wave_all(520) <= 0; 
        tb_wave_all(521) <= 0; 
        tb_wave_all(522) <= 0; 
        tb_wave_all(523) <= 0; 
        tb_wave_all(524) <= 0; 
        tb_wave_all(525) <= 0; 
        tb_wave_all(526) <= 0; 
        tb_wave_all(527) <= 0; 
        tb_wave_all(528) <= 0; 
        tb_wave_all(529) <= 0; 
        tb_wave_all(530) <= 0; 
        tb_wave_all(531) <= 0; 
        tb_wave_all(532) <= 0; 
        tb_wave_all(533) <= 0; 
        tb_wave_all(534) <= 0; 
        tb_wave_all(535) <= 0; 
        tb_wave_all(536) <= 0; 
        tb_wave_all(537) <= 0; 
        tb_wave_all(538) <= 0; 
        tb_wave_all(539) <= 0; 
        tb_wave_all(540) <= 0; 
        tb_wave_all(541) <= 0; 
        tb_wave_all(542) <= 0; 
        tb_wave_all(543) <= 0; 
        tb_wave_all(544) <= 2318; 
        tb_wave_all(545) <= 2685; 
        tb_wave_all(546) <= 2099; 
        tb_wave_all(547) <= 2912; 
        tb_wave_all(548) <= 3756; 
        tb_wave_all(549) <= 3193; 
        tb_wave_all(550) <= 2139; 
        tb_wave_all(551) <= 2335; 
        tb_wave_all(552) <= 0; 
        tb_wave_all(553) <= 0; 
        tb_wave_all(554) <= 0; 
        tb_wave_all(555) <= 0; 
        tb_wave_all(556) <= 0; 
        tb_wave_all(557) <= 0; 
        tb_wave_all(558) <= 0; 
        tb_wave_all(559) <= 0; 
        tb_wave_all(560) <= 0; 
        tb_wave_all(561) <= 0; 
        tb_wave_all(562) <= 0; 
        tb_wave_all(563) <= 0; 
        tb_wave_all(564) <= 0; 
        tb_wave_all(565) <= 0; 
        tb_wave_all(566) <= 0; 
        tb_wave_all(567) <= 0; 
        tb_wave_all(568) <= 0; 
        tb_wave_all(569) <= 0; 
        tb_wave_all(570) <= 0; 
        tb_wave_all(571) <= 0; 
        tb_wave_all(572) <= 0; 
        tb_wave_all(573) <= 0; 
        tb_wave_all(574) <= 0; 
        tb_wave_all(575) <= 0; 
        tb_wave_all(576) <= 64337; 
        tb_wave_all(577) <= 63685; 
        tb_wave_all(578) <= 64143; 
        tb_wave_all(579) <= 64260; 
        tb_wave_all(580) <= 63187; 
        tb_wave_all(581) <= 63236; 
        tb_wave_all(582) <= 63769; 
        tb_wave_all(583) <= 63895; 
        tb_wave_all(584) <= 0; 
        tb_wave_all(585) <= 0; 
        tb_wave_all(586) <= 0; 
        tb_wave_all(587) <= 0; 
        tb_wave_all(588) <= 0; 
        tb_wave_all(589) <= 0; 
        tb_wave_all(590) <= 0; 
        tb_wave_all(591) <= 0; 
        tb_wave_all(592) <= 0; 
        tb_wave_all(593) <= 0; 
        tb_wave_all(594) <= 0; 
        tb_wave_all(595) <= 0; 
        tb_wave_all(596) <= 0; 
        tb_wave_all(597) <= 0; 
        tb_wave_all(598) <= 0; 
        tb_wave_all(599) <= 0; 
        tb_wave_all(600) <= 0; 
        tb_wave_all(601) <= 0; 
        tb_wave_all(602) <= 0; 
        tb_wave_all(603) <= 0; 
        tb_wave_all(604) <= 0; 
        tb_wave_all(605) <= 0; 
        tb_wave_all(606) <= 0; 
        tb_wave_all(607) <= 0; 
        tb_wave_all(608) <= 512; 
        tb_wave_all(609) <= 76; 
        tb_wave_all(610) <= 64904; 
        tb_wave_all(611) <= 64264; 
        tb_wave_all(612) <= 64658; 
        tb_wave_all(613) <= 64123; 
        tb_wave_all(614) <= 62980; 
        tb_wave_all(615) <= 63372; 
        tb_wave_all(616) <= 0; 
        tb_wave_all(617) <= 0; 
        tb_wave_all(618) <= 0; 
        tb_wave_all(619) <= 0; 
        tb_wave_all(620) <= 0; 
        tb_wave_all(621) <= 0; 
        tb_wave_all(622) <= 0; 
        tb_wave_all(623) <= 0; 
        tb_wave_all(624) <= 0; 
        tb_wave_all(625) <= 0; 
        tb_wave_all(626) <= 0; 
        tb_wave_all(627) <= 0; 
        tb_wave_all(628) <= 0; 
        tb_wave_all(629) <= 0; 
        tb_wave_all(630) <= 0; 
        tb_wave_all(631) <= 0; 
        tb_wave_all(632) <= 0; 
        tb_wave_all(633) <= 0; 
        tb_wave_all(634) <= 0; 
        tb_wave_all(635) <= 0; 
        tb_wave_all(636) <= 0; 
        tb_wave_all(637) <= 0; 
        tb_wave_all(638) <= 0; 
        tb_wave_all(639) <= 0; 
        tb_wave_all(640) <= 505; 
        tb_wave_all(641) <= 626; 
        tb_wave_all(642) <= 175; 
        tb_wave_all(643) <= 65440; 
        tb_wave_all(644) <= 634; 
        tb_wave_all(645) <= 65531; 
        tb_wave_all(646) <= 65329; 
        tb_wave_all(647) <= 397; 
        tb_wave_all(648) <= 0; 
        tb_wave_all(649) <= 0; 
        tb_wave_all(650) <= 0; 
        tb_wave_all(651) <= 0; 
        tb_wave_all(652) <= 0; 
        tb_wave_all(653) <= 0; 
        tb_wave_all(654) <= 0; 
        tb_wave_all(655) <= 0; 
        tb_wave_all(656) <= 0; 
        tb_wave_all(657) <= 0; 
        tb_wave_all(658) <= 0; 
        tb_wave_all(659) <= 0; 
        tb_wave_all(660) <= 0; 
        tb_wave_all(661) <= 0; 
        tb_wave_all(662) <= 0; 
        tb_wave_all(663) <= 0; 
        tb_wave_all(664) <= 0; 
        tb_wave_all(665) <= 0; 
        tb_wave_all(666) <= 0; 
        tb_wave_all(667) <= 0; 
        tb_wave_all(668) <= 0; 
        tb_wave_all(669) <= 0; 
        tb_wave_all(670) <= 0; 
        tb_wave_all(671) <= 0; 
        tb_wave_all(672) <= 427; 
        tb_wave_all(673) <= 154; 
        tb_wave_all(674) <= 65243; 
        tb_wave_all(675) <= 64924; 
        tb_wave_all(676) <= 65079; 
        tb_wave_all(677) <= 64987; 
        tb_wave_all(678) <= 64329; 
        tb_wave_all(679) <= 63539; 
        tb_wave_all(680) <= 0; 
        tb_wave_all(681) <= 0; 
        tb_wave_all(682) <= 0; 
        tb_wave_all(683) <= 0; 
        tb_wave_all(684) <= 0; 
        tb_wave_all(685) <= 0; 
        tb_wave_all(686) <= 0; 
        tb_wave_all(687) <= 0; 
        tb_wave_all(688) <= 0; 
        tb_wave_all(689) <= 0; 
        tb_wave_all(690) <= 0; 
        tb_wave_all(691) <= 0; 
        tb_wave_all(692) <= 0; 
        tb_wave_all(693) <= 0; 
        tb_wave_all(694) <= 0; 
        tb_wave_all(695) <= 0; 
        tb_wave_all(696) <= 0; 
        tb_wave_all(697) <= 0; 
        tb_wave_all(698) <= 0; 
        tb_wave_all(699) <= 0; 
        tb_wave_all(700) <= 0; 
        tb_wave_all(701) <= 0; 
        tb_wave_all(702) <= 0; 
        tb_wave_all(703) <= 0; 
        tb_wave_all(704) <= 64933; 
        tb_wave_all(705) <= 65399; 
        tb_wave_all(706) <= 802; 
        tb_wave_all(707) <= 598; 
        tb_wave_all(708) <= 64722; 
        tb_wave_all(709) <= 64974; 
        tb_wave_all(710) <= 65020; 
        tb_wave_all(711) <= 64237; 
        tb_wave_all(712) <= 0; 
        tb_wave_all(713) <= 0; 
        tb_wave_all(714) <= 0; 
        tb_wave_all(715) <= 0; 
        tb_wave_all(716) <= 0; 
        tb_wave_all(717) <= 0; 
        tb_wave_all(718) <= 0; 
        tb_wave_all(719) <= 0; 
        tb_wave_all(720) <= 0; 
        tb_wave_all(721) <= 0; 
        tb_wave_all(722) <= 0; 
        tb_wave_all(723) <= 0; 
        tb_wave_all(724) <= 0; 
        tb_wave_all(725) <= 0; 
        tb_wave_all(726) <= 0; 
        tb_wave_all(727) <= 0; 
        tb_wave_all(728) <= 0; 
        tb_wave_all(729) <= 0; 
        tb_wave_all(730) <= 0; 
        tb_wave_all(731) <= 0; 
        tb_wave_all(732) <= 0; 
        tb_wave_all(733) <= 0; 
        tb_wave_all(734) <= 0; 
        tb_wave_all(735) <= 0; 
        tb_wave_all(736) <= 337; 
        tb_wave_all(737) <= 100; 
        tb_wave_all(738) <= 285; 
        tb_wave_all(739) <= 522; 
        tb_wave_all(740) <= 591; 
        tb_wave_all(741) <= 707; 
        tb_wave_all(742) <= 705; 
        tb_wave_all(743) <= 563; 
        tb_wave_all(744) <= 0; 
        tb_wave_all(745) <= 0; 
        tb_wave_all(746) <= 0; 
        tb_wave_all(747) <= 0; 
        tb_wave_all(748) <= 0; 
        tb_wave_all(749) <= 0; 
        tb_wave_all(750) <= 0; 
        tb_wave_all(751) <= 0; 
        tb_wave_all(752) <= 0; 
        tb_wave_all(753) <= 0; 
        tb_wave_all(754) <= 0; 
        tb_wave_all(755) <= 0; 
        tb_wave_all(756) <= 0; 
        tb_wave_all(757) <= 0; 
        tb_wave_all(758) <= 0; 
        tb_wave_all(759) <= 0; 
        tb_wave_all(760) <= 0; 
        tb_wave_all(761) <= 0; 
        tb_wave_all(762) <= 0; 
        tb_wave_all(763) <= 0; 
        tb_wave_all(764) <= 0; 
        tb_wave_all(765) <= 0; 
        tb_wave_all(766) <= 0; 
        tb_wave_all(767) <= 0; 
        tb_wave_all(768) <= 1506; 
        tb_wave_all(769) <= 2421; 
        tb_wave_all(770) <= 2360; 
        tb_wave_all(771) <= 2157; 
        tb_wave_all(772) <= 3235; 
        tb_wave_all(773) <= 2556; 
        tb_wave_all(774) <= 2045; 
        tb_wave_all(775) <= 3303; 
        tb_wave_all(776) <= 0; 
        tb_wave_all(777) <= 0; 
        tb_wave_all(778) <= 0; 
        tb_wave_all(779) <= 0; 
        tb_wave_all(780) <= 0; 
        tb_wave_all(781) <= 0; 
        tb_wave_all(782) <= 0; 
        tb_wave_all(783) <= 0; 
        tb_wave_all(784) <= 0; 
        tb_wave_all(785) <= 0; 
        tb_wave_all(786) <= 0; 
        tb_wave_all(787) <= 0; 
        tb_wave_all(788) <= 0; 
        tb_wave_all(789) <= 0; 
        tb_wave_all(790) <= 0; 
        tb_wave_all(791) <= 0; 
        tb_wave_all(792) <= 0; 
        tb_wave_all(793) <= 0; 
        tb_wave_all(794) <= 0; 
        tb_wave_all(795) <= 0; 
        tb_wave_all(796) <= 0; 
        tb_wave_all(797) <= 0; 
        tb_wave_all(798) <= 0; 
        tb_wave_all(799) <= 0; 
        tb_wave_all(800) <= 64827; 
        tb_wave_all(801) <= 64938; 
        tb_wave_all(802) <= 65457; 
        tb_wave_all(803) <= 65172; 
        tb_wave_all(804) <= 63778; 
        tb_wave_all(805) <= 63296; 
        tb_wave_all(806) <= 63781; 
        tb_wave_all(807) <= 63938; 
        tb_wave_all(808) <= 0; 
        tb_wave_all(809) <= 0; 
        tb_wave_all(810) <= 0; 
        tb_wave_all(811) <= 0; 
        tb_wave_all(812) <= 0; 
        tb_wave_all(813) <= 0; 
        tb_wave_all(814) <= 0; 
        tb_wave_all(815) <= 0; 
        tb_wave_all(816) <= 0; 
        tb_wave_all(817) <= 0; 
        tb_wave_all(818) <= 0; 
        tb_wave_all(819) <= 0; 
        tb_wave_all(820) <= 0; 
        tb_wave_all(821) <= 0; 
        tb_wave_all(822) <= 0; 
        tb_wave_all(823) <= 0; 
        tb_wave_all(824) <= 0; 
        tb_wave_all(825) <= 0; 
        tb_wave_all(826) <= 0; 
        tb_wave_all(827) <= 0; 
        tb_wave_all(828) <= 0; 
        tb_wave_all(829) <= 0; 
        tb_wave_all(830) <= 0; 
        tb_wave_all(831) <= 0; 
        tb_wave_all(832) <= 65165; 
        tb_wave_all(833) <= 65481; 
        tb_wave_all(834) <= 162; 
        tb_wave_all(835) <= 300; 
        tb_wave_all(836) <= 73; 
        tb_wave_all(837) <= 140; 
        tb_wave_all(838) <= 120; 
        tb_wave_all(839) <= 323; 
        tb_wave_all(840) <= 0; 
        tb_wave_all(841) <= 0; 
        tb_wave_all(842) <= 0; 
        tb_wave_all(843) <= 0; 
        tb_wave_all(844) <= 0; 
        tb_wave_all(845) <= 0; 
        tb_wave_all(846) <= 0; 
        tb_wave_all(847) <= 0; 
        tb_wave_all(848) <= 0; 
        tb_wave_all(849) <= 0; 
        tb_wave_all(850) <= 0; 
        tb_wave_all(851) <= 0; 
        tb_wave_all(852) <= 0; 
        tb_wave_all(853) <= 0; 
        tb_wave_all(854) <= 0; 
        tb_wave_all(855) <= 0; 
        tb_wave_all(856) <= 0; 
        tb_wave_all(857) <= 0; 
        tb_wave_all(858) <= 0; 
        tb_wave_all(859) <= 0; 
        tb_wave_all(860) <= 0; 
        tb_wave_all(861) <= 0; 
        tb_wave_all(862) <= 0; 
        tb_wave_all(863) <= 0; 
        tb_wave_all(864) <= 1155; 
        tb_wave_all(865) <= 1278; 
        tb_wave_all(866) <= 65260; 
        tb_wave_all(867) <= 64511; 
        tb_wave_all(868) <= 65479; 
        tb_wave_all(869) <= 705; 
        tb_wave_all(870) <= 65512; 
        tb_wave_all(871) <= 65142; 
        tb_wave_all(872) <= 0; 
        tb_wave_all(873) <= 0; 
        tb_wave_all(874) <= 0; 
        tb_wave_all(875) <= 0; 
        tb_wave_all(876) <= 0; 
        tb_wave_all(877) <= 0; 
        tb_wave_all(878) <= 0; 
        tb_wave_all(879) <= 0; 
        tb_wave_all(880) <= 0; 
        tb_wave_all(881) <= 0; 
        tb_wave_all(882) <= 0; 
        tb_wave_all(883) <= 0; 
        tb_wave_all(884) <= 0; 
        tb_wave_all(885) <= 0; 
        tb_wave_all(886) <= 0; 
        tb_wave_all(887) <= 0; 
        tb_wave_all(888) <= 0; 
        tb_wave_all(889) <= 0; 
        tb_wave_all(890) <= 0; 
        tb_wave_all(891) <= 0; 
        tb_wave_all(892) <= 0; 
        tb_wave_all(893) <= 0; 
        tb_wave_all(894) <= 0; 
        tb_wave_all(895) <= 0; 
        tb_wave_all(896) <= 1772; 
        tb_wave_all(897) <= 2444; 
        tb_wave_all(898) <= 2505; 
        tb_wave_all(899) <= 1760; 
        tb_wave_all(900) <= 1429; 
        tb_wave_all(901) <= 1114; 
        tb_wave_all(902) <= 207; 
        tb_wave_all(903) <= 65280; 
        tb_wave_all(904) <= 0; 
        tb_wave_all(905) <= 0; 
        tb_wave_all(906) <= 0; 
        tb_wave_all(907) <= 0; 
        tb_wave_all(908) <= 0; 
        tb_wave_all(909) <= 0; 
        tb_wave_all(910) <= 0; 
        tb_wave_all(911) <= 0; 
        tb_wave_all(912) <= 0; 
        tb_wave_all(913) <= 0; 
        tb_wave_all(914) <= 0; 
        tb_wave_all(915) <= 0; 
        tb_wave_all(916) <= 0; 
        tb_wave_all(917) <= 0; 
        tb_wave_all(918) <= 0; 
        tb_wave_all(919) <= 0; 
        tb_wave_all(920) <= 0; 
        tb_wave_all(921) <= 0; 
        tb_wave_all(922) <= 0; 
        tb_wave_all(923) <= 0; 
        tb_wave_all(924) <= 0; 
        tb_wave_all(925) <= 0; 
        tb_wave_all(926) <= 0; 
        tb_wave_all(927) <= 0; 
        tb_wave_all(928) <= 63708; 
        tb_wave_all(929) <= 63765; 
        tb_wave_all(930) <= 64220; 
        tb_wave_all(931) <= 64265; 
        tb_wave_all(932) <= 64572; 
        tb_wave_all(933) <= 64807; 
        tb_wave_all(934) <= 64688; 
        tb_wave_all(935) <= 64973; 
        tb_wave_all(936) <= 0; 
        tb_wave_all(937) <= 0; 
        tb_wave_all(938) <= 0; 
        tb_wave_all(939) <= 0; 
        tb_wave_all(940) <= 0; 
        tb_wave_all(941) <= 0; 
        tb_wave_all(942) <= 0; 
        tb_wave_all(943) <= 0; 
        tb_wave_all(944) <= 0; 
        tb_wave_all(945) <= 0; 
        tb_wave_all(946) <= 0; 
        tb_wave_all(947) <= 0; 
        tb_wave_all(948) <= 0; 
        tb_wave_all(949) <= 0; 
        tb_wave_all(950) <= 0; 
        tb_wave_all(951) <= 0; 
        tb_wave_all(952) <= 0; 
        tb_wave_all(953) <= 0; 
        tb_wave_all(954) <= 0; 
        tb_wave_all(955) <= 0; 
        tb_wave_all(956) <= 0; 
        tb_wave_all(957) <= 0; 
        tb_wave_all(958) <= 0; 
        tb_wave_all(959) <= 0; 
        tb_wave_all(960) <= 1106; 
        tb_wave_all(961) <= 343; 
        tb_wave_all(962) <= 789; 
        tb_wave_all(963) <= 1510; 
        tb_wave_all(964) <= 353; 
        tb_wave_all(965) <= 65151; 
        tb_wave_all(966) <= 309; 
        tb_wave_all(967) <= 842; 
        tb_wave_all(968) <= 0; 
        tb_wave_all(969) <= 0; 
        tb_wave_all(970) <= 0; 
        tb_wave_all(971) <= 0; 
        tb_wave_all(972) <= 0; 
        tb_wave_all(973) <= 0; 
        tb_wave_all(974) <= 0; 
        tb_wave_all(975) <= 0; 
        tb_wave_all(976) <= 0; 
        tb_wave_all(977) <= 0; 
        tb_wave_all(978) <= 0; 
        tb_wave_all(979) <= 0; 
        tb_wave_all(980) <= 0; 
        tb_wave_all(981) <= 0; 
        tb_wave_all(982) <= 0; 
        tb_wave_all(983) <= 0; 
        tb_wave_all(984) <= 0; 
        tb_wave_all(985) <= 0; 
        tb_wave_all(986) <= 0; 
        tb_wave_all(987) <= 0; 
        tb_wave_all(988) <= 0; 
        tb_wave_all(989) <= 0; 
        tb_wave_all(990) <= 0; 
        tb_wave_all(991) <= 0; 
        tb_wave_all(992) <= 2449; 
        tb_wave_all(993) <= 3851; 
        tb_wave_all(994) <= 3561; 
        tb_wave_all(995) <= 3688; 
        tb_wave_all(996) <= 4138; 
        tb_wave_all(997) <= 3217; 
        tb_wave_all(998) <= 3300; 
        tb_wave_all(999) <= 4341; 
        tb_wave_all(1000) <= 0; 
        tb_wave_all(1001) <= 0; 
        tb_wave_all(1002) <= 0; 
        tb_wave_all(1003) <= 0; 
        tb_wave_all(1004) <= 0; 
        tb_wave_all(1005) <= 0; 
        tb_wave_all(1006) <= 0; 
        tb_wave_all(1007) <= 0; 
        tb_wave_all(1008) <= 0; 
        tb_wave_all(1009) <= 0; 
        tb_wave_all(1010) <= 0; 
        tb_wave_all(1011) <= 0; 
        tb_wave_all(1012) <= 0; 
        tb_wave_all(1013) <= 0; 
        tb_wave_all(1014) <= 0; 
        tb_wave_all(1015) <= 0; 
        tb_wave_all(1016) <= 0; 
        tb_wave_all(1017) <= 0; 
        tb_wave_all(1018) <= 0; 
        tb_wave_all(1019) <= 0; 
        tb_wave_all(1020) <= 0; 
        tb_wave_all(1021) <= 0; 
        tb_wave_all(1022) <= 0; 
        tb_wave_all(1023) <= 0; 

        wait for 100 ns;

    end process;

end architecture;